magic
tech sky130A
timestamp 1725973893
<< nwell >>
rect -671 76 73 238
<< nmos >>
rect -571 -96 -556 30
rect -398 -96 -383 30
rect -225 -96 -210 30
rect 0 0 15 42
<< pmos >>
rect -571 94 -556 220
rect -398 94 -383 220
rect -225 94 -210 220
rect 0 94 15 220
<< ndiff >>
rect -611 20 -571 30
rect -611 -2 -601 20
rect -581 -2 -571 20
rect -611 -22 -571 -2
rect -611 -44 -601 -22
rect -581 -44 -571 -22
rect -611 -64 -571 -44
rect -611 -86 -601 -64
rect -581 -86 -571 -64
rect -611 -96 -571 -86
rect -556 20 -516 30
rect -556 -2 -546 20
rect -526 -2 -516 20
rect -556 -22 -516 -2
rect -556 -44 -546 -22
rect -526 -44 -516 -22
rect -556 -64 -516 -44
rect -556 -86 -546 -64
rect -526 -86 -516 -64
rect -556 -96 -516 -86
rect -438 20 -398 30
rect -438 -2 -428 20
rect -408 -2 -398 20
rect -438 -22 -398 -2
rect -438 -44 -428 -22
rect -408 -44 -398 -22
rect -438 -64 -398 -44
rect -438 -86 -428 -64
rect -408 -86 -398 -64
rect -438 -96 -398 -86
rect -383 20 -343 30
rect -383 -2 -373 20
rect -353 -2 -343 20
rect -383 -22 -343 -2
rect -383 -44 -373 -22
rect -353 -44 -343 -22
rect -383 -64 -343 -44
rect -383 -86 -373 -64
rect -353 -86 -343 -64
rect -383 -96 -343 -86
rect -265 20 -225 30
rect -265 -2 -255 20
rect -235 -2 -225 20
rect -265 -22 -225 -2
rect -265 -44 -255 -22
rect -235 -44 -225 -22
rect -265 -64 -225 -44
rect -265 -86 -255 -64
rect -235 -86 -225 -64
rect -265 -96 -225 -86
rect -210 20 -170 30
rect -210 -2 -200 20
rect -180 -2 -170 20
rect -40 32 0 42
rect -40 10 -30 32
rect -10 10 0 32
rect -40 0 0 10
rect 15 32 55 42
rect 15 10 25 32
rect 45 10 55 32
rect 15 0 55 10
rect -210 -22 -170 -2
rect -210 -44 -200 -22
rect -180 -44 -170 -22
rect -210 -64 -170 -44
rect -210 -86 -200 -64
rect -180 -86 -170 -64
rect -210 -96 -170 -86
<< pdiff >>
rect -611 210 -571 220
rect -611 188 -601 210
rect -581 188 -571 210
rect -611 168 -571 188
rect -611 146 -601 168
rect -581 146 -571 168
rect -611 126 -571 146
rect -611 104 -601 126
rect -581 104 -571 126
rect -611 94 -571 104
rect -556 210 -516 220
rect -556 188 -546 210
rect -526 188 -516 210
rect -556 168 -516 188
rect -556 146 -546 168
rect -526 146 -516 168
rect -556 126 -516 146
rect -556 104 -546 126
rect -526 104 -516 126
rect -556 94 -516 104
rect -438 210 -398 220
rect -438 188 -428 210
rect -408 188 -398 210
rect -438 168 -398 188
rect -438 146 -428 168
rect -408 146 -398 168
rect -438 126 -398 146
rect -438 104 -428 126
rect -408 104 -398 126
rect -438 94 -398 104
rect -383 210 -343 220
rect -383 188 -373 210
rect -353 188 -343 210
rect -383 168 -343 188
rect -383 146 -373 168
rect -353 146 -343 168
rect -383 126 -343 146
rect -383 104 -373 126
rect -353 104 -343 126
rect -383 94 -343 104
rect -265 210 -225 220
rect -265 188 -255 210
rect -235 188 -225 210
rect -265 168 -225 188
rect -265 146 -255 168
rect -235 146 -225 168
rect -265 126 -225 146
rect -265 104 -255 126
rect -235 104 -225 126
rect -265 94 -225 104
rect -210 210 -170 220
rect -210 188 -200 210
rect -180 188 -170 210
rect -210 168 -170 188
rect -210 146 -200 168
rect -180 146 -170 168
rect -210 126 -170 146
rect -210 104 -200 126
rect -180 104 -170 126
rect -210 94 -170 104
rect -40 210 0 220
rect -40 188 -30 210
rect -10 188 0 210
rect -40 168 0 188
rect -40 146 -30 168
rect -10 146 0 168
rect -40 126 0 146
rect -40 104 -30 126
rect -10 104 0 126
rect -40 94 0 104
rect 15 210 55 220
rect 15 188 25 210
rect 45 188 55 210
rect 15 168 55 188
rect 15 146 25 168
rect 45 146 55 168
rect 15 126 55 146
rect 15 104 25 126
rect 45 104 55 126
rect 15 94 55 104
<< ndiffc >>
rect -601 -2 -581 20
rect -601 -44 -581 -22
rect -601 -86 -581 -64
rect -546 -2 -526 20
rect -546 -44 -526 -22
rect -546 -86 -526 -64
rect -428 -2 -408 20
rect -428 -44 -408 -22
rect -428 -86 -408 -64
rect -373 -2 -353 20
rect -373 -44 -353 -22
rect -373 -86 -353 -64
rect -255 -2 -235 20
rect -255 -44 -235 -22
rect -255 -86 -235 -64
rect -200 -2 -180 20
rect -30 10 -10 32
rect 25 10 45 32
rect -200 -44 -180 -22
rect -200 -86 -180 -64
<< pdiffc >>
rect -601 188 -581 210
rect -601 146 -581 168
rect -601 104 -581 126
rect -546 188 -526 210
rect -546 146 -526 168
rect -546 104 -526 126
rect -428 188 -408 210
rect -428 146 -408 168
rect -428 104 -408 126
rect -373 188 -353 210
rect -373 146 -353 168
rect -373 104 -353 126
rect -255 188 -235 210
rect -255 146 -235 168
rect -255 104 -235 126
rect -200 188 -180 210
rect -200 146 -180 168
rect -200 104 -180 126
rect -30 188 -10 210
rect -30 146 -10 168
rect -30 104 -10 126
rect 25 188 45 210
rect 25 146 45 168
rect 25 104 45 126
<< psubdiff >>
rect -653 17 -611 30
rect -653 -1 -640 17
rect -622 -1 -611 17
rect -653 -25 -611 -1
rect -653 -43 -640 -25
rect -622 -43 -611 -25
rect -653 -67 -611 -43
rect -653 -85 -640 -67
rect -622 -85 -611 -67
rect -653 -96 -611 -85
rect -480 17 -438 30
rect -480 -1 -467 17
rect -449 -1 -438 17
rect -480 -25 -438 -1
rect -480 -43 -467 -25
rect -449 -43 -438 -25
rect -480 -67 -438 -43
rect -480 -85 -467 -67
rect -449 -85 -438 -67
rect -480 -96 -438 -85
rect -307 17 -265 30
rect -307 -1 -294 17
rect -276 -1 -265 17
rect -307 -25 -265 -1
rect -307 -43 -294 -25
rect -276 -43 -265 -25
rect -307 -67 -265 -43
rect -307 -85 -294 -67
rect -276 -85 -265 -67
rect -307 -96 -265 -85
rect -82 29 -40 42
rect -82 11 -69 29
rect -51 11 -40 29
rect -82 0 -40 11
<< nsubdiff >>
rect -653 207 -611 220
rect -653 189 -640 207
rect -622 189 -611 207
rect -653 165 -611 189
rect -653 147 -640 165
rect -622 147 -611 165
rect -653 123 -611 147
rect -653 105 -640 123
rect -622 105 -611 123
rect -653 94 -611 105
rect -480 207 -438 220
rect -480 189 -467 207
rect -449 189 -438 207
rect -480 165 -438 189
rect -480 147 -467 165
rect -449 147 -438 165
rect -480 123 -438 147
rect -480 105 -467 123
rect -449 105 -438 123
rect -480 94 -438 105
rect -307 207 -265 220
rect -307 189 -294 207
rect -276 189 -265 207
rect -307 165 -265 189
rect -307 147 -294 165
rect -276 147 -265 165
rect -307 123 -265 147
rect -307 105 -294 123
rect -276 105 -265 123
rect -307 94 -265 105
rect -82 207 -40 220
rect -82 189 -69 207
rect -51 189 -40 207
rect -82 165 -40 189
rect -82 147 -69 165
rect -51 147 -40 165
rect -82 123 -40 147
rect -82 105 -69 123
rect -51 105 -40 123
rect -82 94 -40 105
<< psubdiffcont >>
rect -640 -1 -622 17
rect -640 -43 -622 -25
rect -640 -85 -622 -67
rect -467 -1 -449 17
rect -467 -43 -449 -25
rect -467 -85 -449 -67
rect -294 -1 -276 17
rect -294 -43 -276 -25
rect -294 -85 -276 -67
rect -69 11 -51 29
<< nsubdiffcont >>
rect -640 189 -622 207
rect -640 147 -622 165
rect -640 105 -622 123
rect -467 189 -449 207
rect -467 147 -449 165
rect -467 105 -449 123
rect -294 189 -276 207
rect -294 147 -276 165
rect -294 105 -276 123
rect -69 189 -51 207
rect -69 147 -51 165
rect -69 105 -51 123
<< poly >>
rect -571 220 -556 233
rect -398 220 -383 233
rect -225 220 -210 233
rect 0 220 15 233
rect -571 30 -556 94
rect -398 30 -383 94
rect -225 30 -210 94
rect -129 76 -98 84
rect -129 57 -123 76
rect -106 75 -98 76
rect 0 75 15 94
rect -106 60 15 75
rect -106 57 -98 60
rect -129 49 -98 57
rect 0 42 15 60
rect 0 -13 15 0
rect -571 -160 -556 -96
rect -398 -160 -383 -96
rect -225 -160 -210 -96
rect -580 -168 -547 -160
rect -580 -188 -572 -168
rect -555 -188 -547 -168
rect -580 -195 -547 -188
rect -406 -168 -373 -160
rect -406 -188 -398 -168
rect -381 -188 -373 -168
rect -406 -195 -373 -188
rect -234 -168 -201 -160
rect -234 -188 -226 -168
rect -209 -188 -201 -168
rect -234 -195 -201 -188
<< polycont >>
rect -123 57 -106 76
rect -572 -188 -555 -168
rect -398 -188 -381 -168
rect -226 -188 -209 -168
<< locali >>
rect -671 256 -152 260
rect -671 238 -626 256
rect -609 238 -571 256
rect -554 238 -525 256
rect -508 238 -453 256
rect -436 238 -398 256
rect -381 238 -352 256
rect -335 238 -280 256
rect -263 238 -225 256
rect -208 238 -179 256
rect -162 238 -152 256
rect -671 235 -152 238
rect -100 256 73 260
rect -100 238 -55 256
rect -38 238 0 256
rect 17 238 46 256
rect 63 238 73 256
rect -100 235 73 238
rect -671 234 -611 235
rect -498 234 -438 235
rect -325 234 -265 235
rect -100 234 -40 235
rect -646 218 -611 234
rect -473 218 -438 234
rect -300 218 -265 234
rect -75 218 -40 234
rect -646 210 -576 218
rect -646 207 -601 210
rect -646 189 -640 207
rect -622 189 -601 207
rect -646 188 -601 189
rect -581 188 -576 210
rect -646 168 -576 188
rect -646 165 -601 168
rect -646 147 -640 165
rect -622 147 -601 165
rect -646 146 -601 147
rect -581 146 -576 168
rect -646 126 -576 146
rect -646 123 -601 126
rect -646 105 -640 123
rect -622 105 -601 123
rect -646 104 -601 105
rect -581 104 -576 126
rect -646 96 -576 104
rect -554 210 -518 218
rect -554 188 -546 210
rect -526 188 -518 210
rect -554 168 -518 188
rect -554 146 -546 168
rect -526 146 -518 168
rect -554 126 -518 146
rect -554 104 -546 126
rect -526 104 -518 126
rect -554 96 -518 104
rect -473 210 -403 218
rect -473 207 -428 210
rect -473 189 -467 207
rect -449 189 -428 207
rect -473 188 -428 189
rect -408 188 -403 210
rect -473 168 -403 188
rect -473 165 -428 168
rect -473 147 -467 165
rect -449 147 -428 165
rect -473 146 -428 147
rect -408 146 -403 168
rect -473 126 -403 146
rect -473 123 -428 126
rect -473 105 -467 123
rect -449 105 -428 123
rect -473 104 -428 105
rect -408 104 -403 126
rect -473 96 -403 104
rect -381 210 -345 218
rect -381 188 -373 210
rect -353 188 -345 210
rect -381 168 -345 188
rect -381 146 -373 168
rect -353 146 -345 168
rect -381 126 -345 146
rect -381 104 -373 126
rect -353 104 -345 126
rect -381 96 -345 104
rect -300 210 -230 218
rect -300 207 -255 210
rect -300 189 -294 207
rect -276 189 -255 207
rect -300 188 -255 189
rect -235 188 -230 210
rect -300 168 -230 188
rect -300 165 -255 168
rect -300 147 -294 165
rect -276 147 -255 165
rect -300 146 -255 147
rect -235 146 -230 168
rect -300 126 -230 146
rect -300 123 -255 126
rect -300 105 -294 123
rect -276 105 -255 123
rect -300 104 -255 105
rect -235 104 -230 126
rect -300 96 -230 104
rect -208 210 -172 218
rect -208 188 -200 210
rect -180 188 -172 210
rect -208 168 -172 188
rect -208 146 -200 168
rect -180 146 -172 168
rect -208 126 -172 146
rect -208 104 -200 126
rect -180 104 -172 126
rect -208 96 -172 104
rect -75 210 -5 218
rect -75 207 -30 210
rect -75 189 -69 207
rect -51 189 -30 207
rect -75 188 -30 189
rect -10 188 -5 210
rect -75 168 -5 188
rect -75 165 -30 168
rect -75 147 -69 165
rect -51 147 -30 165
rect -75 146 -30 147
rect -10 146 -5 168
rect -75 126 -5 146
rect -75 123 -30 126
rect -75 105 -69 123
rect -51 105 -30 123
rect -75 104 -30 105
rect -10 104 -5 126
rect -75 96 -5 104
rect 17 210 53 218
rect 17 188 25 210
rect 45 188 53 210
rect 17 168 53 188
rect 17 146 25 168
rect 45 146 53 168
rect 17 126 53 146
rect 17 104 25 126
rect 45 104 53 126
rect 17 96 53 104
rect -541 78 -518 96
rect -368 78 -345 96
rect -195 78 -172 96
rect -129 78 -98 84
rect -541 76 -98 78
rect -541 57 -123 76
rect -106 57 -98 76
rect -541 51 -98 57
rect -646 28 -611 30
rect -473 28 -438 30
rect -300 28 -265 30
rect -646 20 -576 28
rect -646 17 -601 20
rect -646 -1 -640 17
rect -622 -1 -601 17
rect -646 -2 -601 -1
rect -581 -2 -576 20
rect -646 -22 -576 -2
rect -646 -25 -601 -22
rect -646 -43 -640 -25
rect -622 -43 -601 -25
rect -646 -44 -601 -43
rect -581 -44 -576 -22
rect -646 -64 -576 -44
rect -646 -67 -601 -64
rect -646 -85 -640 -67
rect -622 -85 -601 -67
rect -646 -86 -601 -85
rect -581 -86 -576 -64
rect -646 -94 -576 -86
rect -554 20 -518 28
rect -554 -2 -546 20
rect -526 -2 -518 20
rect -554 -22 -518 -2
rect -554 -44 -546 -22
rect -526 -44 -518 -22
rect -554 -64 -518 -44
rect -554 -86 -546 -64
rect -526 -79 -518 -64
rect -473 20 -403 28
rect -473 17 -428 20
rect -473 -1 -467 17
rect -449 -1 -428 17
rect -473 -2 -428 -1
rect -408 -2 -403 20
rect -473 -22 -403 -2
rect -473 -25 -428 -22
rect -473 -43 -467 -25
rect -449 -43 -428 -25
rect -473 -44 -428 -43
rect -408 -44 -403 -22
rect -473 -64 -403 -44
rect -473 -67 -428 -64
rect -473 -79 -467 -67
rect -526 -85 -467 -79
rect -449 -85 -428 -67
rect -526 -86 -428 -85
rect -408 -86 -403 -64
rect -554 -94 -403 -86
rect -381 20 -345 28
rect -381 -2 -373 20
rect -353 -2 -345 20
rect -381 -22 -345 -2
rect -381 -44 -373 -22
rect -353 -44 -345 -22
rect -381 -64 -345 -44
rect -381 -86 -373 -64
rect -353 -79 -345 -64
rect -300 20 -230 28
rect -300 17 -255 20
rect -300 -1 -294 17
rect -276 -1 -255 17
rect -300 -2 -255 -1
rect -235 -2 -230 20
rect -300 -22 -230 -2
rect -300 -25 -255 -22
rect -300 -43 -294 -25
rect -276 -43 -255 -25
rect -300 -44 -255 -43
rect -235 -44 -230 -22
rect -300 -64 -230 -44
rect -300 -67 -255 -64
rect -300 -79 -294 -67
rect -353 -85 -294 -79
rect -276 -85 -255 -67
rect -353 -86 -255 -85
rect -235 -86 -230 -64
rect -381 -94 -230 -86
rect -208 20 -172 51
rect -129 49 -98 51
rect 30 40 53 96
rect -208 -2 -200 20
rect -180 -2 -172 20
rect -208 -22 -172 -2
rect -208 -44 -200 -22
rect -180 -44 -172 -22
rect -75 32 -5 40
rect -75 29 -30 32
rect -75 11 -69 29
rect -51 11 -30 29
rect -75 10 -30 11
rect -10 10 -5 32
rect -75 2 -5 10
rect 17 32 53 40
rect 17 10 25 32
rect 45 10 53 32
rect 17 2 53 10
rect -75 -15 -40 2
rect -75 -16 72 -15
rect -75 -34 -55 -16
rect -38 -34 0 -16
rect 17 -34 46 -16
rect 63 -34 72 -16
rect -75 -40 72 -34
rect -208 -64 -172 -44
rect -208 -86 -200 -64
rect -180 -86 -172 -64
rect -208 -94 -172 -86
rect -646 -115 -611 -94
rect -541 -96 -438 -94
rect -368 -96 -265 -94
rect -195 -96 -172 -94
rect -646 -132 -636 -115
rect -619 -132 -607 -115
rect -646 -138 -607 -132
rect -580 -168 -547 -160
rect -580 -188 -572 -168
rect -555 -188 -547 -168
rect -580 -195 -547 -188
rect -406 -168 -373 -160
rect -406 -188 -398 -168
rect -381 -188 -373 -168
rect -406 -195 -373 -188
rect -234 -168 -201 -160
rect -234 -188 -226 -168
rect -209 -188 -201 -168
rect -234 -195 -201 -188
<< viali >>
rect -626 238 -609 256
rect -571 238 -554 256
rect -525 238 -508 256
rect -453 238 -436 256
rect -398 238 -381 256
rect -352 238 -335 256
rect -280 238 -263 256
rect -225 238 -208 256
rect -179 238 -162 256
rect -55 238 -38 256
rect 0 238 17 256
rect 46 238 63 256
rect -55 -34 -38 -16
rect 0 -34 17 -16
rect 46 -34 63 -16
rect -636 -132 -619 -115
<< metal1 >>
rect -671 256 73 260
rect -671 238 -626 256
rect -609 238 -571 256
rect -554 238 -525 256
rect -508 238 -453 256
rect -436 238 -398 256
rect -381 238 -352 256
rect -335 238 -280 256
rect -263 238 -225 256
rect -208 238 -179 256
rect -162 238 -55 256
rect -38 238 0 256
rect 17 238 46 256
rect 63 238 73 256
rect -671 234 73 238
rect -100 -16 73 -13
rect -100 -34 -55 -16
rect -38 -34 0 -16
rect 17 -34 46 -16
rect 63 -34 73 -16
rect -100 -40 73 -34
rect -646 -115 -611 -112
rect -100 -115 -73 -40
rect -646 -132 -636 -115
rect -619 -132 -73 -115
rect -646 -138 -73 -132
<< labels >>
rlabel locali 53 68 53 68 1 y
port 4 n
rlabel locali -218 -192 -218 -192 1 c
port 3 n
rlabel locali -391 -191 -391 -191 1 b
port 2 n
rlabel locali -564 -191 -564 -191 1 a
port 1 n
rlabel metal1 -668 247 -668 247 3 vdd
port 5 e
rlabel metal1 -642 -125 -642 -125 1 vss
port 6 n
<< end >>
