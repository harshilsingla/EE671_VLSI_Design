magic
tech sky130A
timestamp 1726146073
<< nwell >>
rect -1162 142 74 231
<< nmos >>
rect -1064 30 -1049 72
rect -931 30 -916 72
rect -798 30 -783 72
rect -665 30 -650 72
rect -532 30 -517 72
rect -399 30 -384 72
rect -266 30 -251 72
rect -133 30 -118 72
rect 0 30 15 72
<< pmos >>
rect -1064 160 -1049 202
rect -931 160 -916 202
rect -798 160 -783 202
rect -665 160 -650 202
rect -532 160 -517 202
rect -399 160 -384 202
rect -266 160 -251 202
rect -133 160 -118 202
rect 0 160 15 202
<< ndiff >>
rect -1104 61 -1064 72
rect -1104 44 -1094 61
rect -1075 44 -1064 61
rect -1104 30 -1064 44
rect -1049 62 -1009 72
rect -1049 40 -1039 62
rect -1019 40 -1009 62
rect -1049 30 -1009 40
rect -971 62 -931 72
rect -971 40 -961 62
rect -941 40 -931 62
rect -971 30 -931 40
rect -916 62 -876 72
rect -916 40 -906 62
rect -886 40 -876 62
rect -916 30 -876 40
rect -838 62 -798 72
rect -838 40 -828 62
rect -808 40 -798 62
rect -838 30 -798 40
rect -783 62 -743 72
rect -783 40 -773 62
rect -753 40 -743 62
rect -783 30 -743 40
rect -705 62 -665 72
rect -705 40 -695 62
rect -675 40 -665 62
rect -705 30 -665 40
rect -650 62 -610 72
rect -650 40 -640 62
rect -620 40 -610 62
rect -650 30 -610 40
rect -572 62 -532 72
rect -572 40 -562 62
rect -542 40 -532 62
rect -572 30 -532 40
rect -517 62 -477 72
rect -517 40 -507 62
rect -487 40 -477 62
rect -517 30 -477 40
rect -439 61 -399 72
rect -439 44 -430 61
rect -411 44 -399 61
rect -439 30 -399 44
rect -384 62 -344 72
rect -384 45 -374 62
rect -354 45 -344 62
rect -384 30 -344 45
rect -306 62 -266 72
rect -306 45 -297 62
rect -277 45 -266 62
rect -306 30 -266 45
rect -251 63 -211 72
rect -251 46 -241 63
rect -221 46 -211 63
rect -251 30 -211 46
rect -173 62 -133 72
rect -173 40 -163 62
rect -143 40 -133 62
rect -173 30 -133 40
rect -118 62 -78 72
rect -118 40 -108 62
rect -88 40 -78 62
rect -118 30 -78 40
rect -40 62 0 72
rect -40 40 -30 62
rect -10 40 0 62
rect -40 30 0 40
rect 15 62 55 72
rect 15 40 25 62
rect 45 40 55 62
rect 15 30 55 40
<< pdiff >>
rect -1104 192 -1064 202
rect -1104 170 -1094 192
rect -1074 170 -1064 192
rect -1104 160 -1064 170
rect -1049 192 -1009 202
rect -1049 170 -1039 192
rect -1019 170 -1009 192
rect -1049 160 -1009 170
rect -971 192 -931 202
rect -971 170 -961 192
rect -941 170 -931 192
rect -971 160 -931 170
rect -916 192 -876 202
rect -916 170 -906 192
rect -886 170 -876 192
rect -916 160 -876 170
rect -838 192 -798 202
rect -838 170 -828 192
rect -808 170 -798 192
rect -838 160 -798 170
rect -783 192 -743 202
rect -783 170 -773 192
rect -753 170 -743 192
rect -783 160 -743 170
rect -705 192 -665 202
rect -705 170 -695 192
rect -675 170 -665 192
rect -705 160 -665 170
rect -650 192 -610 202
rect -650 170 -640 192
rect -620 170 -610 192
rect -650 160 -610 170
rect -572 192 -532 202
rect -572 170 -562 192
rect -542 170 -532 192
rect -572 160 -532 170
rect -517 192 -477 202
rect -517 170 -507 192
rect -487 170 -477 192
rect -517 160 -477 170
rect -439 192 -399 202
rect -439 170 -429 192
rect -409 170 -399 192
rect -439 160 -399 170
rect -384 192 -344 202
rect -384 170 -374 192
rect -354 170 -344 192
rect -384 160 -344 170
rect -306 192 -266 202
rect -306 170 -296 192
rect -276 170 -266 192
rect -306 160 -266 170
rect -251 192 -211 202
rect -251 170 -241 192
rect -221 170 -211 192
rect -251 160 -211 170
rect -173 192 -133 202
rect -173 170 -163 192
rect -143 170 -133 192
rect -173 160 -133 170
rect -118 192 -78 202
rect -118 170 -108 192
rect -88 170 -78 192
rect -118 160 -78 170
rect -40 192 0 202
rect -40 170 -30 192
rect -10 170 0 192
rect -40 160 0 170
rect 15 192 55 202
rect 15 170 25 192
rect 45 170 55 192
rect 15 160 55 170
<< ndiffc >>
rect -1094 44 -1075 61
rect -1039 40 -1019 62
rect -961 40 -941 62
rect -906 40 -886 62
rect -828 40 -808 62
rect -773 40 -753 62
rect -695 40 -675 62
rect -640 40 -620 62
rect -562 40 -542 62
rect -507 40 -487 62
rect -430 44 -411 61
rect -374 45 -354 62
rect -297 45 -277 62
rect -241 46 -221 63
rect -163 40 -143 62
rect -108 40 -88 62
rect -30 40 -10 62
rect 25 40 45 62
<< pdiffc >>
rect -1094 170 -1074 192
rect -1039 170 -1019 192
rect -961 170 -941 192
rect -906 170 -886 192
rect -828 170 -808 192
rect -773 170 -753 192
rect -695 170 -675 192
rect -640 170 -620 192
rect -562 170 -542 192
rect -507 170 -487 192
rect -429 170 -409 192
rect -374 170 -354 192
rect -296 170 -276 192
rect -241 170 -221 192
rect -163 170 -143 192
rect -108 170 -88 192
rect -30 170 -10 192
rect 25 170 45 192
<< psubdiff >>
rect -1144 60 -1104 72
rect -1144 43 -1132 60
rect -1115 43 -1104 60
rect -1144 30 -1104 43
<< nsubdiff >>
rect -1144 190 -1104 202
rect -1144 170 -1132 190
rect -1115 170 -1104 190
rect -1144 160 -1104 170
<< psubdiffcont >>
rect -1132 43 -1115 60
<< nsubdiffcont >>
rect -1132 170 -1115 190
<< poly >>
rect -1064 202 -1049 218
rect -931 202 -916 218
rect -798 202 -783 218
rect -665 202 -650 218
rect -532 202 -517 218
rect -399 202 -384 218
rect -266 202 -251 218
rect -133 202 -118 218
rect 0 202 15 218
rect -1064 143 -1049 160
rect -931 143 -916 160
rect -798 143 -783 160
rect -1064 128 -783 143
rect -1064 72 -1049 128
rect -931 72 -916 128
rect -798 72 -783 128
rect -665 143 -650 160
rect -532 143 -517 160
rect -399 143 -384 160
rect -665 128 -384 143
rect -665 72 -650 128
rect -532 72 -517 128
rect -399 72 -384 128
rect -266 143 -251 160
rect -133 143 -118 160
rect 0 143 15 160
rect -266 128 15 143
rect -266 72 -251 128
rect -133 72 -118 128
rect 0 72 15 128
rect -1064 16 -1049 30
rect -931 17 -916 30
rect -798 17 -783 30
rect -665 17 -650 30
rect -532 17 -517 30
rect -399 16 -384 30
rect -266 16 -251 30
rect -133 17 -118 30
rect 0 17 15 30
rect -1074 11 -1039 16
rect -1074 -6 -1065 11
rect -1048 -6 -1039 11
rect -1074 -11 -1039 -6
rect -408 11 -373 16
rect -408 -6 -399 11
rect -382 -6 -373 11
rect -408 -11 -373 -6
rect -275 11 -240 16
rect -275 -6 -266 11
rect -249 -6 -240 11
rect -275 -11 -240 -6
<< polycont >>
rect -1065 -6 -1048 11
rect -399 -6 -382 11
rect -266 -6 -249 11
<< locali >>
rect -1123 256 74 259
rect -1123 238 -1064 256
rect -1047 238 -931 256
rect -914 238 -798 256
rect -781 238 -665 256
rect -648 238 -532 256
rect -515 238 -399 256
rect -382 238 -266 256
rect -249 238 -133 256
rect -116 238 0 256
rect 17 238 74 256
rect -1123 235 74 238
rect -1098 200 -1081 235
rect -903 200 -886 235
rect -638 200 -621 235
rect -372 200 -355 235
rect -106 200 -89 235
rect -1102 198 -1069 200
rect -1140 192 -1069 198
rect -1140 190 -1094 192
rect -1140 170 -1132 190
rect -1115 170 -1094 190
rect -1074 170 -1069 192
rect -1140 162 -1069 170
rect -1047 192 -1011 200
rect -1047 170 -1039 192
rect -1019 189 -1011 192
rect -969 192 -936 200
rect -969 189 -961 192
rect -1019 172 -961 189
rect -1019 170 -1011 172
rect -1047 162 -1011 170
rect -969 170 -961 172
rect -941 170 -936 192
rect -969 162 -936 170
rect -914 192 -878 200
rect -914 170 -906 192
rect -886 188 -878 192
rect -836 192 -803 200
rect -836 188 -828 192
rect -886 171 -828 188
rect -886 170 -878 171
rect -914 162 -878 170
rect -836 170 -828 171
rect -808 170 -803 192
rect -836 162 -803 170
rect -781 192 -745 200
rect -781 170 -773 192
rect -753 189 -745 192
rect -703 192 -670 200
rect -703 189 -695 192
rect -753 172 -695 189
rect -753 170 -745 172
rect -781 162 -745 170
rect -703 170 -695 172
rect -675 170 -670 192
rect -703 162 -670 170
rect -648 192 -612 200
rect -648 170 -640 192
rect -620 190 -612 192
rect -570 192 -537 200
rect -570 190 -562 192
rect -620 173 -562 190
rect -620 170 -612 173
rect -648 162 -612 170
rect -570 170 -562 173
rect -542 170 -537 192
rect -570 162 -537 170
rect -515 192 -479 200
rect -515 170 -507 192
rect -487 189 -479 192
rect -437 192 -404 200
rect -437 189 -429 192
rect -487 172 -429 189
rect -487 170 -479 172
rect -515 162 -479 170
rect -437 170 -429 172
rect -409 170 -404 192
rect -437 162 -404 170
rect -382 192 -346 200
rect -382 170 -374 192
rect -354 189 -346 192
rect -304 192 -271 200
rect -304 189 -296 192
rect -354 172 -296 189
rect -354 170 -346 172
rect -382 162 -346 170
rect -304 170 -296 172
rect -276 170 -271 192
rect -304 162 -271 170
rect -249 192 -213 200
rect -249 170 -241 192
rect -221 188 -213 192
rect -171 192 -138 200
rect -171 188 -163 192
rect -221 171 -163 188
rect -221 170 -213 171
rect -249 162 -213 170
rect -171 170 -163 171
rect -143 170 -138 192
rect -171 162 -138 170
rect -116 192 -80 200
rect -116 170 -108 192
rect -88 189 -80 192
rect -38 192 -5 200
rect -38 189 -30 192
rect -88 172 -30 189
rect -88 170 -80 172
rect -116 162 -80 170
rect -38 170 -30 172
rect -10 170 -5 192
rect -38 162 -5 170
rect 17 192 53 200
rect 17 170 25 192
rect 45 170 53 192
rect 17 162 53 170
rect -1094 144 -1073 145
rect -1094 127 -1092 144
rect -1075 127 -1073 144
rect -1094 125 -1073 127
rect -1038 144 -1021 162
rect -1092 70 -1075 125
rect -1038 124 -1021 127
rect -903 70 -886 145
rect -771 144 -754 162
rect -771 124 -754 127
rect -505 144 -488 162
rect -505 124 -488 127
rect -239 144 -222 162
rect -239 125 -222 127
rect 27 144 44 162
rect 27 126 44 127
rect -560 87 -88 104
rect -560 70 -543 87
rect -105 70 -88 87
rect -1102 67 -1069 70
rect -1140 61 -1069 67
rect -1140 60 -1094 61
rect -1140 43 -1132 60
rect -1115 44 -1094 60
rect -1075 44 -1069 61
rect -1115 43 -1069 44
rect -1140 35 -1069 43
rect -1102 34 -1069 35
rect -1047 62 -1011 70
rect -1047 40 -1039 62
rect -1019 51 -1011 62
rect -969 62 -936 70
rect -969 51 -961 62
rect -1019 40 -961 51
rect -941 40 -936 62
rect -1047 34 -936 40
rect -1016 32 -936 34
rect -914 62 -878 70
rect -914 40 -906 62
rect -886 58 -878 62
rect -836 62 -803 70
rect -836 58 -828 62
rect -886 41 -828 58
rect -886 40 -878 41
rect -914 32 -878 40
rect -836 40 -828 41
rect -808 40 -803 62
rect -836 32 -803 40
rect -781 62 -745 70
rect -781 40 -773 62
rect -753 57 -745 62
rect -703 62 -670 70
rect -703 57 -695 62
rect -753 40 -695 57
rect -675 40 -670 62
rect -781 32 -745 40
rect -703 32 -670 40
rect -648 62 -612 70
rect -648 40 -640 62
rect -620 59 -612 62
rect -570 62 -537 70
rect -570 59 -562 62
rect -620 42 -562 59
rect -620 40 -612 42
rect -648 32 -612 40
rect -570 40 -562 42
rect -542 40 -537 62
rect -570 32 -537 40
rect -515 62 -479 70
rect -515 40 -507 62
rect -487 53 -479 62
rect -437 61 -404 70
rect -437 53 -430 61
rect -487 44 -430 53
rect -411 44 -404 61
rect -487 40 -404 44
rect -515 35 -404 40
rect -382 62 -346 70
rect -382 45 -374 62
rect -354 61 -346 62
rect -304 62 -271 70
rect -304 61 -297 62
rect -354 45 -297 61
rect -277 45 -271 62
rect -382 44 -271 45
rect -382 35 -346 44
rect -515 34 -421 35
rect -515 32 -425 34
rect -304 33 -271 44
rect -249 63 -213 70
rect -249 46 -241 63
rect -221 60 -213 63
rect -171 62 -138 70
rect -171 60 -163 62
rect -221 46 -163 60
rect -249 43 -163 46
rect -249 33 -213 43
rect -171 40 -163 43
rect -143 40 -138 62
rect -171 32 -138 40
rect -116 62 -80 70
rect -116 40 -108 62
rect -88 59 -80 62
rect -38 62 -5 70
rect -38 59 -30 62
rect -88 42 -30 59
rect -88 40 -80 42
rect -116 32 -80 40
rect -38 40 -30 42
rect -10 40 -5 62
rect -38 32 -5 40
rect 17 62 53 70
rect 17 40 25 62
rect 45 40 53 62
rect 17 32 53 40
rect -1074 11 -1039 16
rect -1074 -6 -1065 11
rect -1048 -6 -1039 11
rect -1001 15 -984 32
rect -467 15 -450 32
rect -1001 -2 -450 15
rect -408 11 -373 16
rect -1074 -11 -1039 -6
rect -408 -6 -399 11
rect -382 -6 -373 11
rect -408 -11 -373 -6
rect -275 11 -240 16
rect -275 -6 -266 11
rect -249 -6 -240 11
rect -275 -11 -240 -6
rect -162 -13 -145 32
rect 27 -13 44 32
rect -207 -16 74 -13
rect -207 -34 -133 -16
rect -116 -34 0 -16
rect 17 -34 74 -16
rect -207 -37 74 -34
<< viali >>
rect -1064 238 -1047 256
rect -931 238 -914 256
rect -798 238 -781 256
rect -665 238 -648 256
rect -532 238 -515 256
rect -399 238 -382 256
rect -266 238 -249 256
rect -133 238 -116 256
rect 0 238 17 256
rect -1092 127 -1075 144
rect -1038 127 -1021 144
rect -771 127 -754 144
rect -505 127 -488 144
rect -239 127 -222 144
rect 27 127 44 144
rect -133 -34 -116 -16
rect 0 -34 17 -16
<< metal1 >>
rect -1123 256 74 259
rect -1123 238 -1064 256
rect -1047 238 -931 256
rect -914 238 -798 256
rect -781 238 -665 256
rect -648 238 -532 256
rect -515 238 -399 256
rect -382 238 -266 256
rect -249 238 -133 256
rect -116 238 0 256
rect 17 238 74 256
rect -1123 235 74 238
rect -1125 144 72 147
rect -1125 127 -1092 144
rect -1075 127 -1038 144
rect -1021 127 -771 144
rect -754 127 -505 144
rect -488 127 -239 144
rect -222 127 27 144
rect 44 127 72 144
rect -1125 123 72 127
rect -1123 -16 74 -13
rect -1123 -34 -133 -16
rect -116 -34 0 -16
rect 17 -34 74 -16
rect -1123 -37 74 -34
<< labels >>
rlabel polycont -1056 2 -1056 2 1 a
port 1 n
rlabel polycont -391 1 -391 1 1 b
port 2 n
rlabel polycont -258 2 -258 2 1 c
port 3 n
rlabel metal1 62 135 62 135 1 y
port 4 n
rlabel metal1 55 247 55 247 1 vdd
port 5 n
rlabel metal1 59 -27 59 -27 1 vss
port 6 n
<< end >>
