* NGSPICE file created from and3.ext - technology: sky130A

.subckt and3 a b c y vdd vss
X0 vdd b y vdd sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.64 as=0.186667 ps=1.822222 w=0.42 l=0.15
**devattr s=1680,164 d=1680,164
X1 a_n1049_30# a y y sky130_fd_pr__nfet_01v8 ad=0.168 pd=1.64 as=0.168 ps=1.64 w=0.42 l=0.15
**devattr s=1680,164 d=1680,164
X2 vdd a y vdd sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.64 as=0.186667 ps=1.822222 w=0.42 l=0.15
**devattr s=1680,164 d=1680,164
X3 y c vdd vdd sky130_fd_pr__pfet_01v8 ad=0.186667 pd=1.822222 as=0.168 ps=1.64 w=0.42 l=0.15
**devattr s=1680,164 d=1680,164
X4 y c vdd vdd sky130_fd_pr__pfet_01v8 ad=0.186667 pd=1.822222 as=0.168 ps=1.64 w=0.42 l=0.15
**devattr s=1680,164 d=1680,164
X5 vss c a_n650_30# y sky130_fd_pr__nfet_01v8 ad=0.168 pd=1.64 as=0.168 ps=1.64 w=0.42 l=0.15
**devattr s=1680,164 d=1680,164
X6 a_n916_30# a a_n1049_30# y sky130_fd_pr__nfet_01v8 ad=0.168 pd=1.64 as=0.168 ps=1.64 w=0.42 l=0.15
**devattr s=1680,164 d=1680,164
X7 a_n1049_30# b a_n650_30# y sky130_fd_pr__nfet_01v8 ad=0.168 pd=1.64 as=0.168 ps=1.64 w=0.42 l=0.15
**devattr s=1680,164 d=1680,164
X8 a_n650_30# c vss y sky130_fd_pr__nfet_01v8 ad=0.168 pd=1.64 as=0.168 ps=1.64 w=0.42 l=0.15
**devattr s=1680,164 d=1680,164
X9 y a vdd vdd sky130_fd_pr__pfet_01v8 ad=0.186667 pd=1.822222 as=0.168 ps=1.64 w=0.42 l=0.15
**devattr s=1680,164 d=1680,164
X10 y b vdd vdd sky130_fd_pr__pfet_01v8 ad=0.186667 pd=1.822222 as=0.168 ps=1.64 w=0.42 l=0.15
**devattr s=1680,164 d=1680,164
X11 y a vdd vdd sky130_fd_pr__pfet_01v8 ad=0.186667 pd=1.822222 as=0.168 ps=1.64 w=0.42 l=0.15
**devattr s=1680,164 d=1680,164
X12 a_n650_30# b a_n783_30# y sky130_fd_pr__nfet_01v8 ad=0.168 pd=1.64 as=0.168 ps=1.64 w=0.42 l=0.15
**devattr s=1680,164 d=1680,164
X13 vss c a_n384_30# y sky130_fd_pr__nfet_01v8 ad=0.168 pd=1.64 as=0.168 ps=1.64 w=0.42 l=0.15
**devattr s=1680,164 d=1680,164
X14 a_n783_30# a a_n916_30# y sky130_fd_pr__nfet_01v8 ad=0.168 pd=1.64 as=0.168 ps=1.64 w=0.42 l=0.15
**devattr s=1680,164 d=1680,164
X15 a_n384_30# b a_n1049_30# y sky130_fd_pr__nfet_01v8 ad=0.168 pd=1.64 as=0.168 ps=1.64 w=0.42 l=0.15
**devattr s=1680,164 d=1680,164
X16 vdd b y vdd sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.64 as=0.186667 ps=1.822222 w=0.42 l=0.15
**devattr s=1680,164 d=1680,164
X17 vdd c y vdd sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.64 as=0.186667 ps=1.822222 w=0.42 l=0.15
**devattr s=1680,164 d=1680,164
.ends

