magic
tech sky130A
timestamp 1726119572
<< nwell >>
rect -564 238 -300 239
rect -721 76 73 238
rect -564 74 -300 76
<< nmos >>
rect -621 -96 -606 30
rect -423 -96 -408 30
rect -225 -96 -210 30
rect 0 0 15 42
<< pmos >>
rect -621 94 -606 220
rect -423 94 -408 220
rect -225 94 -210 220
rect 0 94 15 220
<< ndiff >>
rect -40 32 0 42
rect -661 20 -621 30
rect -661 -2 -651 20
rect -631 -2 -621 20
rect -661 -22 -621 -2
rect -661 -44 -651 -22
rect -631 -44 -621 -22
rect -661 -64 -621 -44
rect -661 -86 -651 -64
rect -631 -86 -621 -64
rect -661 -96 -621 -86
rect -606 20 -566 30
rect -606 -2 -596 20
rect -576 -2 -566 20
rect -606 -22 -566 -2
rect -606 -44 -596 -22
rect -576 -44 -566 -22
rect -606 -64 -566 -44
rect -606 -86 -596 -64
rect -576 -86 -566 -64
rect -606 -96 -566 -86
rect -463 20 -423 30
rect -463 -2 -453 20
rect -433 -2 -423 20
rect -463 -22 -423 -2
rect -463 -44 -453 -22
rect -433 -44 -423 -22
rect -463 -64 -423 -44
rect -463 -86 -453 -64
rect -433 -86 -423 -64
rect -463 -96 -423 -86
rect -408 20 -368 30
rect -408 -2 -398 20
rect -378 -2 -368 20
rect -408 -22 -368 -2
rect -408 -44 -398 -22
rect -378 -44 -368 -22
rect -408 -64 -368 -44
rect -408 -86 -398 -64
rect -378 -86 -368 -64
rect -408 -96 -368 -86
rect -265 20 -225 30
rect -265 -2 -255 20
rect -235 -2 -225 20
rect -265 -22 -225 -2
rect -265 -44 -255 -22
rect -235 -44 -225 -22
rect -265 -64 -225 -44
rect -265 -86 -255 -64
rect -235 -86 -225 -64
rect -265 -96 -225 -86
rect -210 20 -170 30
rect -210 -2 -200 20
rect -180 -2 -170 20
rect -40 10 -30 32
rect -10 10 0 32
rect -40 0 0 10
rect 15 32 55 42
rect 15 10 25 32
rect 45 10 55 32
rect 15 0 55 10
rect -210 -22 -170 -2
rect -210 -44 -200 -22
rect -180 -44 -170 -22
rect -210 -64 -170 -44
rect -210 -86 -200 -64
rect -180 -86 -170 -64
rect -210 -96 -170 -86
<< pdiff >>
rect -661 210 -621 220
rect -661 188 -651 210
rect -631 188 -621 210
rect -661 168 -621 188
rect -661 146 -651 168
rect -631 146 -621 168
rect -661 126 -621 146
rect -661 104 -651 126
rect -631 104 -621 126
rect -661 94 -621 104
rect -606 210 -566 220
rect -606 188 -596 210
rect -576 188 -566 210
rect -606 168 -566 188
rect -606 146 -596 168
rect -576 146 -566 168
rect -606 126 -566 146
rect -606 104 -596 126
rect -576 104 -566 126
rect -606 94 -566 104
rect -463 210 -423 220
rect -463 188 -453 210
rect -433 188 -423 210
rect -463 168 -423 188
rect -463 146 -453 168
rect -433 146 -423 168
rect -463 126 -423 146
rect -463 104 -453 126
rect -433 104 -423 126
rect -463 94 -423 104
rect -408 210 -368 220
rect -408 188 -398 210
rect -378 188 -368 210
rect -408 168 -368 188
rect -408 146 -398 168
rect -378 146 -368 168
rect -408 126 -368 146
rect -408 104 -398 126
rect -378 104 -368 126
rect -408 94 -368 104
rect -265 210 -225 220
rect -265 188 -255 210
rect -235 188 -225 210
rect -265 168 -225 188
rect -265 146 -255 168
rect -235 146 -225 168
rect -265 126 -225 146
rect -265 104 -255 126
rect -235 104 -225 126
rect -265 94 -225 104
rect -210 210 -170 220
rect -210 188 -200 210
rect -180 188 -170 210
rect -210 168 -170 188
rect -210 146 -200 168
rect -180 146 -170 168
rect -210 126 -170 146
rect -210 104 -200 126
rect -180 104 -170 126
rect -210 94 -170 104
rect -40 210 0 220
rect -40 188 -30 210
rect -10 188 0 210
rect -40 168 0 188
rect -40 146 -30 168
rect -10 146 0 168
rect -40 126 0 146
rect -40 104 -30 126
rect -10 104 0 126
rect -40 94 0 104
rect 15 210 55 220
rect 15 188 25 210
rect 45 188 55 210
rect 15 168 55 188
rect 15 146 25 168
rect 45 146 55 168
rect 15 126 55 146
rect 15 104 25 126
rect 45 104 55 126
rect 15 94 55 104
<< ndiffc >>
rect -651 -2 -631 20
rect -651 -44 -631 -22
rect -651 -86 -631 -64
rect -596 -2 -576 20
rect -596 -44 -576 -22
rect -596 -86 -576 -64
rect -453 -2 -433 20
rect -453 -44 -433 -22
rect -453 -86 -433 -64
rect -398 -2 -378 20
rect -398 -44 -378 -22
rect -398 -86 -378 -64
rect -255 -2 -235 20
rect -255 -44 -235 -22
rect -255 -86 -235 -64
rect -200 -2 -180 20
rect -30 10 -10 32
rect 25 10 45 32
rect -200 -44 -180 -22
rect -200 -86 -180 -64
<< pdiffc >>
rect -651 188 -631 210
rect -651 146 -631 168
rect -651 104 -631 126
rect -596 188 -576 210
rect -596 146 -576 168
rect -596 104 -576 126
rect -453 188 -433 210
rect -453 146 -433 168
rect -453 104 -433 126
rect -398 188 -378 210
rect -398 146 -378 168
rect -398 104 -378 126
rect -255 188 -235 210
rect -255 146 -235 168
rect -255 104 -235 126
rect -200 188 -180 210
rect -200 146 -180 168
rect -200 104 -180 126
rect -30 188 -10 210
rect -30 146 -10 168
rect -30 104 -10 126
rect 25 188 45 210
rect 25 146 45 168
rect 25 104 45 126
<< psubdiff >>
rect -703 17 -661 30
rect -703 -1 -690 17
rect -672 -1 -661 17
rect -703 -25 -661 -1
rect -703 -43 -690 -25
rect -672 -43 -661 -25
rect -703 -67 -661 -43
rect -703 -85 -690 -67
rect -672 -85 -661 -67
rect -703 -96 -661 -85
<< nsubdiff >>
rect -703 207 -661 220
rect -703 189 -690 207
rect -672 189 -661 207
rect -703 165 -661 189
rect -703 147 -690 165
rect -672 147 -661 165
rect -703 123 -661 147
rect -703 105 -690 123
rect -672 105 -661 123
rect -703 94 -661 105
<< psubdiffcont >>
rect -690 -1 -672 17
rect -690 -43 -672 -25
rect -690 -85 -672 -67
<< nsubdiffcont >>
rect -690 189 -672 207
rect -690 147 -672 165
rect -690 105 -672 123
<< poly >>
rect -621 220 -606 233
rect -423 220 -408 233
rect -225 220 -210 233
rect 0 220 15 233
rect -621 30 -606 94
rect -423 30 -408 94
rect -225 30 -210 94
rect -129 76 -98 84
rect -129 57 -123 76
rect -106 75 -98 76
rect 0 75 15 94
rect -106 60 15 75
rect -106 57 -98 60
rect -129 49 -98 57
rect 0 42 15 60
rect 0 -13 15 0
rect -621 -160 -606 -96
rect -423 -160 -408 -96
rect -225 -160 -210 -96
rect -630 -168 -597 -160
rect -630 -188 -622 -168
rect -605 -188 -597 -168
rect -630 -195 -597 -188
rect -431 -168 -398 -160
rect -431 -188 -423 -168
rect -406 -188 -398 -168
rect -431 -195 -398 -188
rect -234 -168 -201 -160
rect -234 -188 -226 -168
rect -209 -188 -201 -168
rect -234 -195 -201 -188
<< polycont >>
rect -123 57 -106 76
rect -622 -188 -605 -168
rect -423 -188 -406 -168
rect -226 -188 -209 -168
<< locali >>
rect -721 256 -152 260
rect -721 238 -676 256
rect -659 238 -621 256
rect -604 238 -575 256
rect -558 238 -478 256
rect -461 238 -423 256
rect -406 238 -377 256
rect -360 238 -280 256
rect -263 238 -225 256
rect -208 238 -179 256
rect -162 238 -152 256
rect -721 237 -152 238
rect -721 235 -379 237
rect -352 235 -152 237
rect -100 256 73 260
rect -100 238 -55 256
rect -38 238 0 256
rect 17 238 46 256
rect 63 238 73 256
rect -100 235 73 238
rect -721 234 -661 235
rect -548 234 -463 235
rect -352 234 -265 235
rect -100 234 -40 235
rect -696 218 -661 234
rect -498 218 -463 234
rect -300 218 -265 234
rect -75 218 -40 234
rect -696 210 -626 218
rect -696 207 -651 210
rect -696 189 -690 207
rect -672 189 -651 207
rect -696 188 -651 189
rect -631 188 -626 210
rect -696 168 -626 188
rect -696 165 -651 168
rect -696 147 -690 165
rect -672 147 -651 165
rect -696 146 -651 147
rect -631 146 -626 168
rect -696 126 -626 146
rect -696 123 -651 126
rect -696 105 -690 123
rect -672 105 -651 123
rect -696 104 -651 105
rect -631 104 -626 126
rect -696 96 -626 104
rect -604 210 -568 218
rect -604 188 -596 210
rect -576 188 -568 210
rect -604 168 -568 188
rect -604 146 -596 168
rect -576 146 -568 168
rect -604 126 -568 146
rect -604 104 -596 126
rect -576 104 -568 126
rect -604 96 -568 104
rect -498 210 -428 218
rect -498 188 -453 210
rect -433 188 -428 210
rect -498 168 -428 188
rect -498 146 -453 168
rect -433 146 -428 168
rect -498 126 -428 146
rect -498 104 -453 126
rect -433 104 -428 126
rect -498 96 -428 104
rect -406 210 -370 218
rect -406 188 -398 210
rect -378 188 -370 210
rect -406 168 -370 188
rect -406 146 -398 168
rect -378 146 -370 168
rect -406 126 -370 146
rect -406 104 -398 126
rect -378 104 -370 126
rect -406 96 -370 104
rect -300 210 -230 218
rect -300 188 -255 210
rect -235 188 -230 210
rect -300 168 -230 188
rect -300 146 -255 168
rect -235 146 -230 168
rect -300 126 -230 146
rect -300 104 -255 126
rect -235 104 -230 126
rect -300 96 -230 104
rect -208 210 -172 218
rect -208 188 -200 210
rect -180 188 -172 210
rect -208 168 -172 188
rect -208 146 -200 168
rect -180 146 -172 168
rect -208 126 -172 146
rect -208 104 -200 126
rect -180 104 -172 126
rect -208 96 -172 104
rect -75 210 -5 218
rect -75 188 -30 210
rect -10 188 -5 210
rect -75 168 -5 188
rect -75 146 -30 168
rect -10 146 -5 168
rect -75 126 -5 146
rect -75 104 -30 126
rect -10 104 -5 126
rect -75 96 -5 104
rect 17 210 53 218
rect 17 188 25 210
rect 45 188 53 210
rect 17 168 53 188
rect 17 146 25 168
rect 45 146 53 168
rect 17 126 53 146
rect 17 104 25 126
rect 45 104 53 126
rect 17 96 53 104
rect -591 78 -568 96
rect -393 78 -370 96
rect -195 78 -172 96
rect -129 78 -98 84
rect -591 77 -542 78
rect -517 77 -349 78
rect -324 77 -98 78
rect -591 76 -98 77
rect -591 57 -123 76
rect -106 57 -98 76
rect -591 51 -98 57
rect -552 49 -511 51
rect -357 49 -316 51
rect -696 28 -661 30
rect -498 28 -463 30
rect -300 28 -265 30
rect -696 20 -626 28
rect -696 17 -651 20
rect -696 -1 -690 17
rect -672 -1 -651 17
rect -696 -2 -651 -1
rect -631 -2 -626 20
rect -696 -22 -626 -2
rect -696 -25 -651 -22
rect -696 -43 -690 -25
rect -672 -43 -651 -25
rect -696 -44 -651 -43
rect -631 -44 -626 -22
rect -696 -64 -626 -44
rect -696 -67 -651 -64
rect -696 -85 -690 -67
rect -672 -85 -651 -67
rect -696 -86 -651 -85
rect -631 -86 -626 -64
rect -696 -94 -626 -86
rect -604 20 -568 28
rect -604 -2 -596 20
rect -576 -2 -568 20
rect -604 -22 -568 -2
rect -604 -44 -596 -22
rect -576 -44 -568 -22
rect -604 -64 -568 -44
rect -604 -86 -596 -64
rect -576 -72 -568 -64
rect -498 20 -428 28
rect -498 -2 -453 20
rect -433 -2 -428 20
rect -498 -22 -428 -2
rect -498 -44 -453 -22
rect -433 -44 -428 -22
rect -498 -64 -428 -44
rect -498 -71 -453 -64
rect -576 -78 -544 -72
rect -576 -86 -564 -78
rect -604 -94 -564 -86
rect -696 -115 -661 -94
rect -591 -95 -564 -94
rect -547 -95 -544 -78
rect -591 -96 -544 -95
rect -570 -101 -544 -96
rect -527 -77 -453 -71
rect -527 -94 -523 -77
rect -506 -86 -453 -77
rect -433 -86 -428 -64
rect -506 -94 -428 -86
rect -406 20 -370 28
rect -406 -2 -398 20
rect -378 -2 -370 20
rect -406 -22 -370 -2
rect -406 -44 -398 -22
rect -378 -44 -370 -22
rect -406 -64 -370 -44
rect -300 20 -230 28
rect -300 -2 -255 20
rect -235 -2 -230 20
rect -300 -22 -230 -2
rect -300 -44 -255 -22
rect -235 -44 -230 -22
rect -300 -64 -230 -44
rect -406 -86 -398 -64
rect -378 -75 -343 -64
rect -300 -68 -255 -64
rect -378 -86 -368 -75
rect -406 -92 -368 -86
rect -351 -90 -343 -75
rect -326 -77 -255 -68
rect -351 -92 -344 -90
rect -406 -94 -344 -92
rect -527 -96 -463 -94
rect -393 -96 -344 -94
rect -326 -94 -322 -77
rect -305 -86 -255 -77
rect -235 -86 -230 -64
rect -305 -94 -230 -86
rect -208 20 -172 51
rect -129 49 -98 51
rect 30 40 53 96
rect -208 -2 -200 20
rect -180 -2 -172 20
rect -208 -22 -172 -2
rect -208 -44 -200 -22
rect -180 -44 -172 -22
rect -75 32 -5 40
rect -75 10 -30 32
rect -10 10 -5 32
rect -75 2 -5 10
rect 17 32 53 40
rect 17 10 25 32
rect 45 10 53 32
rect 17 2 53 10
rect -75 -15 -40 2
rect -75 -16 72 -15
rect -75 -34 -55 -16
rect -38 -34 0 -16
rect 17 -34 46 -16
rect 63 -34 72 -16
rect -75 -40 72 -34
rect -208 -64 -172 -44
rect -208 -86 -200 -64
rect -180 -86 -172 -64
rect -208 -94 -172 -86
rect -326 -96 -265 -94
rect -195 -96 -172 -94
rect -527 -100 -501 -96
rect -326 -101 -294 -96
rect -696 -132 -686 -115
rect -669 -132 -657 -115
rect -696 -138 -657 -132
rect -630 -168 -597 -160
rect -630 -188 -622 -168
rect -605 -188 -597 -168
rect -630 -195 -597 -188
rect -431 -168 -398 -160
rect -431 -188 -423 -168
rect -406 -188 -398 -168
rect -431 -195 -398 -188
rect -234 -168 -201 -160
rect -234 -188 -226 -168
rect -209 -188 -201 -168
rect -234 -195 -201 -188
<< viali >>
rect -676 238 -659 256
rect -621 238 -604 256
rect -575 238 -558 256
rect -478 238 -461 256
rect -423 238 -406 256
rect -377 238 -360 256
rect -280 238 -263 256
rect -225 238 -208 256
rect -179 238 -162 256
rect -55 238 -38 256
rect 0 238 17 256
rect 46 238 63 256
rect -564 -95 -547 -78
rect -523 -94 -506 -77
rect -368 -92 -351 -75
rect -322 -94 -305 -77
rect -55 -34 -38 -16
rect 0 -34 17 -16
rect 46 -34 63 -16
rect -686 -132 -669 -115
<< metal1 >>
rect -721 256 73 260
rect -721 238 -676 256
rect -659 238 -621 256
rect -604 238 -575 256
rect -558 238 -478 256
rect -461 238 -423 256
rect -406 238 -377 256
rect -360 238 -280 256
rect -263 238 -225 256
rect -208 238 -179 256
rect -162 238 -55 256
rect -38 238 0 256
rect 17 238 46 256
rect 63 238 73 256
rect -721 234 73 238
rect -100 -16 73 -13
rect -100 -34 -55 -16
rect -38 -34 0 -16
rect 17 -34 46 -16
rect 63 -34 73 -16
rect -100 -40 73 -34
rect -375 -68 -343 -64
rect -570 -78 -544 -72
rect -570 -95 -564 -78
rect -547 -79 -544 -78
rect -527 -77 -501 -71
rect -527 -79 -523 -77
rect -547 -94 -523 -79
rect -506 -94 -501 -77
rect -547 -95 -501 -94
rect -570 -96 -501 -95
rect -375 -75 -294 -68
rect -375 -92 -368 -75
rect -351 -77 -294 -75
rect -351 -92 -322 -77
rect -375 -94 -322 -92
rect -305 -94 -294 -77
rect -375 -96 -294 -94
rect -570 -101 -544 -96
rect -527 -100 -501 -96
rect -357 -99 -294 -96
rect -326 -101 -294 -99
rect -696 -115 -661 -112
rect -100 -115 -73 -40
rect -696 -132 -686 -115
rect -669 -132 -73 -115
rect -696 -138 -73 -132
<< labels >>
rlabel locali 53 68 53 68 1 y
port 4 n
rlabel locali -218 -192 -218 -192 1 c
port 3 n
rlabel locali -614 -191 -614 -191 1 a
port 1 n
rlabel metal1 -718 247 -718 247 3 vdd
port 5 e
rlabel metal1 -692 -125 -692 -125 1 vss
port 6 n
rlabel locali -416 -191 -416 -191 1 b
port 2 n
rlabel viali -553 -89 -553 -89 1 temp1
port 7 n
rlabel viali -356 -86 -356 -86 1 temp2
port 8 n
<< end >>
