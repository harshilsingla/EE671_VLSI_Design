magic
tech sky130A
timestamp 1726158675
<< nwell >>
rect -100 76 73 238
<< nmos >>
rect 0 0 15 42
<< pmos >>
rect 0 94 15 220
<< ndiff >>
rect -40 32 0 42
rect -40 10 -30 32
rect -10 10 0 32
rect -40 0 0 10
rect 15 32 55 42
rect 15 10 25 32
rect 45 10 55 32
rect 15 0 55 10
<< pdiff >>
rect -40 210 0 220
rect -40 188 -30 210
rect -10 188 0 210
rect -40 168 0 188
rect -40 146 -30 168
rect -10 146 0 168
rect -40 126 0 146
rect -40 104 -30 126
rect -10 104 0 126
rect -40 94 0 104
rect 15 210 55 220
rect 15 188 25 210
rect 45 188 55 210
rect 15 168 55 188
rect 15 146 25 168
rect 45 146 55 168
rect 15 126 55 146
rect 15 104 25 126
rect 45 104 55 126
rect 15 94 55 104
<< ndiffc >>
rect -30 10 -10 32
rect 25 10 45 32
<< pdiffc >>
rect -30 188 -10 210
rect -30 146 -10 168
rect -30 104 -10 126
rect 25 188 45 210
rect 25 146 45 168
rect 25 104 45 126
<< psubdiff >>
rect -82 29 -40 42
rect -82 11 -69 29
rect -51 11 -40 29
rect -82 0 -40 11
<< nsubdiff >>
rect -82 207 -40 220
rect -82 189 -69 207
rect -51 189 -40 207
rect -82 165 -40 189
rect -82 147 -69 165
rect -51 147 -40 165
rect -82 123 -40 147
rect -82 105 -69 123
rect -51 105 -40 123
rect -82 94 -40 105
<< psubdiffcont >>
rect -69 11 -51 29
<< nsubdiffcont >>
rect -69 189 -51 207
rect -69 147 -51 165
rect -69 105 -51 123
<< poly >>
rect 0 220 15 233
rect -129 76 -98 84
rect -129 57 -123 76
rect -106 75 -98 76
rect 0 75 15 94
rect -106 60 15 75
rect -106 57 -98 60
rect -129 49 -98 57
rect 0 42 15 60
rect 0 -13 15 0
<< polycont >>
rect -123 57 -106 76
<< locali >>
rect -100 256 73 259
rect -100 238 -55 256
rect -38 238 0 256
rect 17 238 46 256
rect 63 238 73 256
rect -100 235 73 238
rect -100 234 -40 235
rect -75 218 -40 234
rect -75 210 -5 218
rect -75 207 -30 210
rect -75 189 -69 207
rect -51 189 -30 207
rect -75 188 -30 189
rect -10 188 -5 210
rect -75 168 -5 188
rect -75 165 -30 168
rect -75 147 -69 165
rect -51 147 -30 165
rect -75 146 -30 147
rect -10 146 -5 168
rect -75 126 -5 146
rect -75 123 -30 126
rect -75 105 -69 123
rect -51 105 -30 123
rect -75 104 -30 105
rect -10 104 -5 126
rect -75 96 -5 104
rect 17 210 53 218
rect 17 188 25 210
rect 45 188 53 210
rect 17 168 53 188
rect 17 146 25 168
rect 45 146 53 168
rect 17 126 53 146
rect 17 104 25 126
rect 45 104 53 126
rect 17 96 53 104
rect -129 76 -98 84
rect -129 57 -123 76
rect -106 57 -98 76
rect -129 49 -98 57
rect 30 40 53 96
rect -75 32 -5 40
rect -75 29 -30 32
rect -75 11 -69 29
rect -51 11 -30 29
rect -75 10 -30 11
rect -10 10 -5 32
rect -75 2 -5 10
rect 17 32 53 40
rect 17 10 25 32
rect 45 10 53 32
rect 17 2 53 10
rect -75 -13 -40 2
rect -100 -15 -40 -13
rect -100 -16 72 -15
rect -100 -34 -55 -16
rect -38 -34 0 -16
rect 17 -34 46 -16
rect 63 -34 72 -16
rect -100 -37 72 -34
<< viali >>
rect -55 238 -38 256
rect 0 238 17 256
rect 46 238 63 256
rect -55 -34 -38 -16
rect 0 -34 17 -16
rect 46 -34 63 -16
<< metal1 >>
rect -100 256 73 259
rect -100 238 -55 256
rect -38 238 0 256
rect 17 238 46 256
rect 63 238 73 256
rect -100 234 73 238
rect -100 -16 73 -13
rect -100 -34 -55 -16
rect -38 -34 0 -16
rect 17 -34 46 -16
rect 63 -34 73 -16
rect -100 -37 73 -34
<< labels >>
rlabel metal1 -100 247 -100 247 1 vdd
port 2 n
rlabel metal1 -100 -26 -100 -26 1 vss
port 1 n
rlabel locali -123 67 -123 67 1 a
port 3 n
rlabel locali 53 68 53 68 1 y
port 4 n
<< end >>
