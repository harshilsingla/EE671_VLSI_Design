* NGSPICE file created from inverter.ext - technology: sky130A

X0 y a vss vss sky130_fd_pr__nfet_01v8 ad=0.168 pd=1.64 as=0.168 ps=1.64 w=0.42 l=0.15
X1 y a vdd vdd sky130_fd_pr__pfet_01v8 ad=0.504 pd=3.32 as=0.504 ps=3.32 w=1.26 l=0.15
C0 a vdd 0.119273f
C1 a y 0.031239f
C2 y vdd 0.146586f
C3 y vss 0.168883f
C4 a vss 0.333831f
C5 vdd vss 0.633345f
