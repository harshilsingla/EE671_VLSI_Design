* SkyWater PDK

.subckt inverter vss vdd a y
xm01  y a  vdd vdd sky130_fd_pr__pfet_01v8 l=0.15 w=1.26 
xm02  y a  vss vss sky130_fd_pr__nfet_01v8 l=0.15 w=0.42 
.ends

.subckt inv2 vss vdd a y
Xinverter_0 vss vdd a y inverter
Xinverter_1 vss vdd a y inverter
.ends
