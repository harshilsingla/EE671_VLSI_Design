magic
tech sky130A
timestamp 1726158675
<< nwell >>
rect -1112 137 157 226
<< nmos >>
rect -1014 25 -999 67
rect -881 25 -866 67
rect -748 25 -733 67
rect -615 25 -600 67
rect -482 25 -467 67
rect -349 25 -334 67
rect -216 25 -201 67
rect -83 25 -68 67
rect 50 25 65 67
<< pmos >>
rect -1014 155 -999 197
rect -881 155 -866 197
rect -748 155 -733 197
rect -615 155 -600 197
rect -482 155 -467 197
rect -349 155 -334 197
rect -216 155 -201 197
rect -83 155 -68 197
rect 50 155 65 197
<< ndiff >>
rect -1054 56 -1014 67
rect -1054 39 -1044 56
rect -1025 39 -1014 56
rect -1054 25 -1014 39
rect -999 57 -959 67
rect -999 35 -989 57
rect -969 35 -959 57
rect -999 25 -959 35
rect -921 57 -881 67
rect -921 35 -911 57
rect -891 35 -881 57
rect -921 25 -881 35
rect -866 57 -826 67
rect -866 35 -856 57
rect -836 35 -826 57
rect -866 25 -826 35
rect -788 57 -748 67
rect -788 35 -778 57
rect -758 35 -748 57
rect -788 25 -748 35
rect -733 57 -693 67
rect -733 35 -723 57
rect -703 35 -693 57
rect -733 25 -693 35
rect -655 57 -615 67
rect -655 35 -645 57
rect -625 35 -615 57
rect -655 25 -615 35
rect -600 57 -560 67
rect -600 35 -590 57
rect -570 35 -560 57
rect -600 25 -560 35
rect -522 57 -482 67
rect -522 35 -512 57
rect -492 35 -482 57
rect -522 25 -482 35
rect -467 57 -427 67
rect -467 35 -457 57
rect -437 35 -427 57
rect -467 25 -427 35
rect -389 56 -349 67
rect -389 39 -380 56
rect -361 39 -349 56
rect -389 25 -349 39
rect -334 57 -294 67
rect -334 40 -324 57
rect -304 40 -294 57
rect -334 25 -294 40
rect -256 57 -216 67
rect -256 40 -247 57
rect -227 40 -216 57
rect -256 25 -216 40
rect -201 58 -161 67
rect -201 41 -191 58
rect -171 41 -161 58
rect -201 25 -161 41
rect -123 57 -83 67
rect -123 35 -113 57
rect -93 35 -83 57
rect -123 25 -83 35
rect -68 57 -28 67
rect -68 35 -58 57
rect -38 35 -28 57
rect -68 25 -28 35
rect 10 57 50 67
rect 10 35 20 57
rect 40 35 50 57
rect 10 25 50 35
rect 65 57 105 67
rect 65 35 75 57
rect 95 35 105 57
rect 65 25 105 35
<< pdiff >>
rect -1054 187 -1014 197
rect -1054 165 -1044 187
rect -1024 165 -1014 187
rect -1054 155 -1014 165
rect -999 187 -959 197
rect -999 165 -989 187
rect -969 165 -959 187
rect -999 155 -959 165
rect -921 187 -881 197
rect -921 165 -911 187
rect -891 165 -881 187
rect -921 155 -881 165
rect -866 187 -826 197
rect -866 165 -856 187
rect -836 165 -826 187
rect -866 155 -826 165
rect -788 187 -748 197
rect -788 165 -778 187
rect -758 165 -748 187
rect -788 155 -748 165
rect -733 187 -693 197
rect -733 165 -723 187
rect -703 165 -693 187
rect -733 155 -693 165
rect -655 187 -615 197
rect -655 165 -645 187
rect -625 165 -615 187
rect -655 155 -615 165
rect -600 187 -560 197
rect -600 165 -590 187
rect -570 165 -560 187
rect -600 155 -560 165
rect -522 187 -482 197
rect -522 165 -512 187
rect -492 165 -482 187
rect -522 155 -482 165
rect -467 187 -427 197
rect -467 165 -457 187
rect -437 165 -427 187
rect -467 155 -427 165
rect -389 187 -349 197
rect -389 165 -379 187
rect -359 165 -349 187
rect -389 155 -349 165
rect -334 187 -294 197
rect -334 165 -324 187
rect -304 165 -294 187
rect -334 155 -294 165
rect -256 187 -216 197
rect -256 165 -246 187
rect -226 165 -216 187
rect -256 155 -216 165
rect -201 187 -161 197
rect -201 165 -191 187
rect -171 165 -161 187
rect -201 155 -161 165
rect -123 187 -83 197
rect -123 165 -113 187
rect -93 165 -83 187
rect -123 155 -83 165
rect -68 187 -28 197
rect -68 165 -58 187
rect -38 165 -28 187
rect -68 155 -28 165
rect 10 187 50 197
rect 10 165 20 187
rect 40 165 50 187
rect 10 155 50 165
rect 65 187 105 197
rect 65 165 75 187
rect 95 165 105 187
rect 65 155 105 165
<< ndiffc >>
rect -1044 39 -1025 56
rect -989 35 -969 57
rect -911 35 -891 57
rect -856 35 -836 57
rect -778 35 -758 57
rect -723 35 -703 57
rect -645 35 -625 57
rect -590 35 -570 57
rect -512 35 -492 57
rect -457 35 -437 57
rect -380 39 -361 56
rect -324 40 -304 57
rect -247 40 -227 57
rect -191 41 -171 58
rect -113 35 -93 57
rect -58 35 -38 57
rect 20 35 40 57
rect 75 35 95 57
<< pdiffc >>
rect -1044 165 -1024 187
rect -989 165 -969 187
rect -911 165 -891 187
rect -856 165 -836 187
rect -778 165 -758 187
rect -723 165 -703 187
rect -645 165 -625 187
rect -590 165 -570 187
rect -512 165 -492 187
rect -457 165 -437 187
rect -379 165 -359 187
rect -324 165 -304 187
rect -246 165 -226 187
rect -191 165 -171 187
rect -113 165 -93 187
rect -58 165 -38 187
rect 20 165 40 187
rect 75 165 95 187
<< psubdiff >>
rect -1094 55 -1054 67
rect -1094 38 -1082 55
rect -1065 38 -1054 55
rect -1094 25 -1054 38
<< nsubdiff >>
rect -1094 185 -1054 197
rect -1094 165 -1082 185
rect -1065 165 -1054 185
rect -1094 155 -1054 165
<< psubdiffcont >>
rect -1082 38 -1065 55
<< nsubdiffcont >>
rect -1082 165 -1065 185
<< poly >>
rect -1014 197 -999 213
rect -881 197 -866 213
rect -748 197 -733 213
rect -615 197 -600 213
rect -482 197 -467 213
rect -349 197 -334 213
rect -216 197 -201 213
rect -83 197 -68 213
rect 50 197 65 213
rect -1014 138 -999 155
rect -881 138 -866 155
rect -748 138 -733 155
rect -1014 123 -733 138
rect -1014 67 -999 123
rect -881 67 -866 123
rect -748 67 -733 123
rect -615 138 -600 155
rect -482 138 -467 155
rect -349 138 -334 155
rect -615 123 -334 138
rect -615 67 -600 123
rect -482 67 -467 123
rect -349 67 -334 123
rect -216 138 -201 155
rect -83 138 -68 155
rect 50 138 65 155
rect -216 123 65 138
rect -216 67 -201 123
rect -83 67 -68 123
rect 50 67 65 123
rect -1014 11 -999 25
rect -881 12 -866 25
rect -748 12 -733 25
rect -615 12 -600 25
rect -482 12 -467 25
rect -349 11 -334 25
rect -216 11 -201 25
rect -83 12 -68 25
rect 50 12 65 25
rect -1024 6 -989 11
rect -1024 -11 -1015 6
rect -998 -11 -989 6
rect -1024 -16 -989 -11
rect -358 6 -323 11
rect -358 -11 -349 6
rect -332 -11 -323 6
rect -358 -16 -323 -11
rect -225 6 -190 11
rect -225 -11 -216 6
rect -199 -11 -190 6
rect -225 -16 -190 -11
<< polycont >>
rect -1015 -11 -998 6
rect -349 -11 -332 6
rect -216 -11 -199 6
<< locali >>
rect -1112 251 151 254
rect -1112 233 -1014 251
rect -997 233 -881 251
rect -864 233 -748 251
rect -731 233 -615 251
rect -598 233 -482 251
rect -465 233 -349 251
rect -332 233 -216 251
rect -199 233 -83 251
rect -66 233 50 251
rect 67 233 151 251
rect -1112 230 151 233
rect -1048 195 -1031 230
rect -853 195 -836 230
rect -588 195 -571 230
rect -322 195 -305 230
rect -56 195 -39 230
rect -1052 193 -1019 195
rect -1090 187 -1019 193
rect -1090 185 -1044 187
rect -1090 165 -1082 185
rect -1065 165 -1044 185
rect -1024 165 -1019 187
rect -1090 157 -1019 165
rect -997 187 -961 195
rect -997 165 -989 187
rect -969 184 -961 187
rect -919 187 -886 195
rect -919 184 -911 187
rect -969 167 -911 184
rect -969 165 -961 167
rect -997 157 -961 165
rect -919 165 -911 167
rect -891 165 -886 187
rect -919 157 -886 165
rect -864 187 -828 195
rect -864 165 -856 187
rect -836 183 -828 187
rect -786 187 -753 195
rect -786 183 -778 187
rect -836 166 -778 183
rect -836 165 -828 166
rect -864 157 -828 165
rect -786 165 -778 166
rect -758 165 -753 187
rect -786 157 -753 165
rect -731 187 -695 195
rect -731 165 -723 187
rect -703 184 -695 187
rect -653 187 -620 195
rect -653 184 -645 187
rect -703 167 -645 184
rect -703 165 -695 167
rect -731 157 -695 165
rect -653 165 -645 167
rect -625 165 -620 187
rect -653 157 -620 165
rect -598 187 -562 195
rect -598 165 -590 187
rect -570 185 -562 187
rect -520 187 -487 195
rect -520 185 -512 187
rect -570 168 -512 185
rect -570 165 -562 168
rect -598 157 -562 165
rect -520 165 -512 168
rect -492 165 -487 187
rect -520 157 -487 165
rect -465 187 -429 195
rect -465 165 -457 187
rect -437 184 -429 187
rect -387 187 -354 195
rect -387 184 -379 187
rect -437 167 -379 184
rect -437 165 -429 167
rect -465 157 -429 165
rect -387 165 -379 167
rect -359 165 -354 187
rect -387 157 -354 165
rect -332 187 -296 195
rect -332 165 -324 187
rect -304 184 -296 187
rect -254 187 -221 195
rect -254 184 -246 187
rect -304 167 -246 184
rect -304 165 -296 167
rect -332 157 -296 165
rect -254 165 -246 167
rect -226 165 -221 187
rect -254 157 -221 165
rect -199 187 -163 195
rect -199 165 -191 187
rect -171 183 -163 187
rect -121 187 -88 195
rect -121 183 -113 187
rect -171 166 -113 183
rect -171 165 -163 166
rect -199 157 -163 165
rect -121 165 -113 166
rect -93 165 -88 187
rect -121 157 -88 165
rect -66 187 -30 195
rect -66 165 -58 187
rect -38 184 -30 187
rect 12 187 45 195
rect 12 184 20 187
rect -38 167 20 184
rect -38 165 -30 167
rect -66 157 -30 165
rect 12 165 20 167
rect 40 165 45 187
rect 12 157 45 165
rect 67 187 103 195
rect 67 165 75 187
rect 95 165 103 187
rect 67 157 103 165
rect -1044 139 -1023 140
rect -1044 122 -1042 139
rect -1025 122 -1023 139
rect -1044 120 -1023 122
rect -988 139 -971 157
rect -1042 65 -1025 120
rect -988 119 -971 122
rect -853 65 -836 140
rect -721 139 -704 157
rect -721 119 -704 122
rect -455 139 -438 157
rect -455 119 -438 122
rect -189 139 -172 157
rect -189 120 -172 122
rect 77 139 94 157
rect 77 121 94 122
rect -510 82 -38 99
rect -510 65 -493 82
rect -55 65 -38 82
rect -1052 62 -1019 65
rect -1090 56 -1019 62
rect -1090 55 -1044 56
rect -1090 38 -1082 55
rect -1065 39 -1044 55
rect -1025 39 -1019 56
rect -1065 38 -1019 39
rect -1090 30 -1019 38
rect -1052 29 -1019 30
rect -997 57 -961 65
rect -997 35 -989 57
rect -969 46 -961 57
rect -919 57 -886 65
rect -919 46 -911 57
rect -969 35 -911 46
rect -891 35 -886 57
rect -997 29 -886 35
rect -966 27 -886 29
rect -864 57 -828 65
rect -864 35 -856 57
rect -836 53 -828 57
rect -786 57 -753 65
rect -786 53 -778 57
rect -836 36 -778 53
rect -836 35 -828 36
rect -864 27 -828 35
rect -786 35 -778 36
rect -758 35 -753 57
rect -786 27 -753 35
rect -731 57 -695 65
rect -731 35 -723 57
rect -703 52 -695 57
rect -653 57 -620 65
rect -653 52 -645 57
rect -703 35 -645 52
rect -625 35 -620 57
rect -731 27 -695 35
rect -653 27 -620 35
rect -598 57 -562 65
rect -598 35 -590 57
rect -570 54 -562 57
rect -520 57 -487 65
rect -520 54 -512 57
rect -570 37 -512 54
rect -570 35 -562 37
rect -598 27 -562 35
rect -520 35 -512 37
rect -492 35 -487 57
rect -520 27 -487 35
rect -465 57 -429 65
rect -465 35 -457 57
rect -437 48 -429 57
rect -387 56 -354 65
rect -387 48 -380 56
rect -437 39 -380 48
rect -361 39 -354 56
rect -437 35 -354 39
rect -465 30 -354 35
rect -332 57 -296 65
rect -332 40 -324 57
rect -304 56 -296 57
rect -254 57 -221 65
rect -254 56 -247 57
rect -304 40 -247 56
rect -227 40 -221 57
rect -332 39 -221 40
rect -332 30 -296 39
rect -465 29 -371 30
rect -465 27 -375 29
rect -254 28 -221 39
rect -199 58 -163 65
rect -199 41 -191 58
rect -171 55 -163 58
rect -121 57 -88 65
rect -121 55 -113 57
rect -171 41 -113 55
rect -199 38 -113 41
rect -199 28 -163 38
rect -121 35 -113 38
rect -93 35 -88 57
rect -121 27 -88 35
rect -66 57 -30 65
rect -66 35 -58 57
rect -38 54 -30 57
rect 12 57 45 65
rect 12 54 20 57
rect -38 37 20 54
rect -38 35 -30 37
rect -66 27 -30 35
rect 12 35 20 37
rect 40 35 45 57
rect 12 27 45 35
rect 67 57 103 65
rect 67 35 75 57
rect 95 35 103 57
rect 67 27 103 35
rect -1024 6 -989 11
rect -1024 -11 -1015 6
rect -998 -11 -989 6
rect -951 10 -934 27
rect -417 10 -400 27
rect -951 -7 -400 10
rect -358 6 -323 11
rect -1024 -16 -989 -11
rect -358 -11 -349 6
rect -332 -11 -323 6
rect -358 -16 -323 -11
rect -225 6 -190 11
rect -225 -11 -216 6
rect -199 -11 -190 6
rect -225 -16 -190 -11
rect -112 -18 -95 27
rect 77 -18 94 27
rect 121 -18 156 -17
rect -157 -21 156 -18
rect -157 -39 -83 -21
rect -66 -39 50 -21
rect 67 -39 156 -21
rect -157 -42 156 -39
<< viali >>
rect -1014 233 -997 251
rect -881 233 -864 251
rect -748 233 -731 251
rect -615 233 -598 251
rect -482 233 -465 251
rect -349 233 -332 251
rect -216 233 -199 251
rect -83 233 -66 251
rect 50 233 67 251
rect -1042 122 -1025 139
rect -988 122 -971 139
rect -721 122 -704 139
rect -455 122 -438 139
rect -189 122 -172 139
rect 77 122 94 139
rect 126 52 143 71
rect -83 -39 -66 -21
rect 50 -39 67 -21
<< metal1 >>
rect -1112 251 151 254
rect -1112 233 -1014 251
rect -997 233 -881 251
rect -864 233 -748 251
rect -731 233 -615 251
rect -598 233 -482 251
rect -465 233 -349 251
rect -332 233 -216 251
rect -199 233 -83 251
rect -66 233 50 251
rect 67 233 151 251
rect -1112 230 151 233
rect -1075 139 141 142
rect -1075 122 -1042 139
rect -1025 122 -988 139
rect -971 122 -721 139
rect -704 122 -455 139
rect -438 122 -189 139
rect -172 122 77 139
rect 94 122 141 139
rect -1075 118 141 122
rect 126 79 141 118
rect 120 71 151 79
rect 120 52 126 71
rect 143 52 151 71
rect 120 45 151 52
rect 121 -18 156 -17
rect -1112 -21 156 -18
rect -1112 -39 -83 -21
rect -66 -39 50 -21
rect 67 -39 156 -21
rect -1112 -42 156 -39
use inverter  inverter_0 ~/Desktop/skywater/Project_1/inv
timestamp 1726158675
transform 1 0 249 0 1 -5
box -129 -37 73 259
<< labels >>
rlabel metal1 109 -32 109 -32 1 vss
port 6 n
rlabel metal1 105 242 105 242 1 vdd
port 5 n
rlabel polycont -208 -3 -208 -3 1 c
port 3 n
rlabel polycont -341 -4 -341 -4 1 b
port 2 n
rlabel polycont -1006 -3 -1006 -3 1 a
port 1 n
rlabel space 292 66 292 66 1 y
port 4 n
<< end >>
