magic
tech sky130A
timestamp 1726347566
<< nwell >>
rect -100 76 583 238
<< nmos >>
rect 0 0 15 42
rect 170 0 185 42
rect 340 0 355 42
rect 510 0 525 42
<< pmos >>
rect 0 94 15 220
rect 170 94 185 220
rect 340 94 355 220
rect 510 94 525 220
<< ndiff >>
rect -40 32 0 42
rect -40 10 -30 32
rect -10 10 0 32
rect -40 0 0 10
rect 15 32 55 42
rect 15 10 25 32
rect 45 10 55 32
rect 15 0 55 10
rect 130 32 170 42
rect 130 10 140 32
rect 160 10 170 32
rect 130 0 170 10
rect 185 32 225 42
rect 185 10 195 32
rect 215 10 225 32
rect 185 0 225 10
rect 300 32 340 42
rect 300 10 310 32
rect 330 10 340 32
rect 300 0 340 10
rect 355 32 395 42
rect 355 10 365 32
rect 385 10 395 32
rect 355 0 395 10
rect 470 32 510 42
rect 470 10 480 32
rect 500 10 510 32
rect 470 0 510 10
rect 525 32 565 42
rect 525 10 535 32
rect 555 10 565 32
rect 525 0 565 10
<< pdiff >>
rect -40 210 0 220
rect -40 188 -30 210
rect -10 188 0 210
rect -40 168 0 188
rect -40 146 -30 168
rect -10 146 0 168
rect -40 126 0 146
rect -40 104 -30 126
rect -10 104 0 126
rect -40 94 0 104
rect 15 210 55 220
rect 15 188 25 210
rect 45 188 55 210
rect 15 168 55 188
rect 15 146 25 168
rect 45 146 55 168
rect 15 126 55 146
rect 15 104 25 126
rect 45 104 55 126
rect 15 94 55 104
rect 130 210 170 220
rect 130 188 140 210
rect 160 188 170 210
rect 130 168 170 188
rect 130 146 140 168
rect 160 146 170 168
rect 130 126 170 146
rect 130 104 140 126
rect 160 104 170 126
rect 130 94 170 104
rect 185 210 225 220
rect 185 188 195 210
rect 215 188 225 210
rect 185 168 225 188
rect 185 146 195 168
rect 215 146 225 168
rect 185 126 225 146
rect 185 104 195 126
rect 215 104 225 126
rect 185 94 225 104
rect 300 210 340 220
rect 300 188 310 210
rect 330 188 340 210
rect 300 168 340 188
rect 300 146 310 168
rect 330 146 340 168
rect 300 126 340 146
rect 300 104 310 126
rect 330 104 340 126
rect 300 94 340 104
rect 355 210 395 220
rect 355 188 365 210
rect 385 188 395 210
rect 355 168 395 188
rect 355 146 365 168
rect 385 146 395 168
rect 355 126 395 146
rect 355 104 365 126
rect 385 104 395 126
rect 355 94 395 104
rect 470 210 510 220
rect 470 188 480 210
rect 500 188 510 210
rect 470 168 510 188
rect 470 146 480 168
rect 500 146 510 168
rect 470 126 510 146
rect 470 104 480 126
rect 500 104 510 126
rect 470 94 510 104
rect 525 210 565 220
rect 525 188 535 210
rect 555 188 565 210
rect 525 168 565 188
rect 525 146 535 168
rect 555 146 565 168
rect 525 126 565 146
rect 525 104 535 126
rect 555 104 565 126
rect 525 94 565 104
<< ndiffc >>
rect -30 10 -10 32
rect 25 10 45 32
rect 140 10 160 32
rect 195 10 215 32
rect 310 10 330 32
rect 365 10 385 32
rect 480 10 500 32
rect 535 10 555 32
<< pdiffc >>
rect -30 188 -10 210
rect -30 146 -10 168
rect -30 104 -10 126
rect 25 188 45 210
rect 25 146 45 168
rect 25 104 45 126
rect 140 188 160 210
rect 140 146 160 168
rect 140 104 160 126
rect 195 188 215 210
rect 195 146 215 168
rect 195 104 215 126
rect 310 188 330 210
rect 310 146 330 168
rect 310 104 330 126
rect 365 188 385 210
rect 365 146 385 168
rect 365 104 385 126
rect 480 188 500 210
rect 480 146 500 168
rect 480 104 500 126
rect 535 188 555 210
rect 535 146 555 168
rect 535 104 555 126
<< psubdiff >>
rect -82 29 -40 42
rect -82 11 -69 29
rect -51 11 -40 29
rect -82 0 -40 11
rect 88 29 130 42
rect 88 11 101 29
rect 119 11 130 29
rect 88 0 130 11
rect 258 29 300 42
rect 258 11 271 29
rect 289 11 300 29
rect 258 0 300 11
rect 428 29 470 42
rect 428 11 441 29
rect 459 11 470 29
rect 428 0 470 11
<< nsubdiff >>
rect -82 207 -40 220
rect -82 189 -69 207
rect -51 189 -40 207
rect -82 165 -40 189
rect -82 147 -69 165
rect -51 147 -40 165
rect -82 123 -40 147
rect -82 105 -69 123
rect -51 105 -40 123
rect -82 94 -40 105
rect 88 207 130 220
rect 88 189 101 207
rect 119 189 130 207
rect 88 165 130 189
rect 88 147 101 165
rect 119 147 130 165
rect 88 123 130 147
rect 88 105 101 123
rect 119 105 130 123
rect 88 94 130 105
rect 258 207 300 220
rect 258 189 271 207
rect 289 189 300 207
rect 258 165 300 189
rect 258 147 271 165
rect 289 147 300 165
rect 258 123 300 147
rect 258 105 271 123
rect 289 105 300 123
rect 258 94 300 105
rect 428 207 470 220
rect 428 189 441 207
rect 459 189 470 207
rect 428 165 470 189
rect 428 147 441 165
rect 459 147 470 165
rect 428 123 470 147
rect 428 105 441 123
rect 459 105 470 123
rect 428 94 470 105
<< psubdiffcont >>
rect -69 11 -51 29
rect 101 11 119 29
rect 271 11 289 29
rect 441 11 459 29
<< nsubdiffcont >>
rect -69 189 -51 207
rect -69 147 -51 165
rect -69 105 -51 123
rect 101 189 119 207
rect 101 147 119 165
rect 101 105 119 123
rect 271 189 289 207
rect 271 147 289 165
rect 271 105 289 123
rect 441 189 459 207
rect 441 147 459 165
rect 441 105 459 123
<< poly >>
rect 0 220 15 233
rect 170 220 185 233
rect 340 220 355 233
rect 510 220 525 233
rect -137 75 -101 83
rect 0 75 15 94
rect 170 75 185 94
rect 340 75 355 94
rect 510 75 525 94
rect -137 55 -129 75
rect -109 60 525 75
rect -109 55 -101 60
rect -137 47 -101 55
rect 0 42 15 60
rect 170 42 185 60
rect 340 42 355 60
rect 510 42 525 60
rect 0 -13 15 0
rect 170 -13 185 0
rect 340 -13 355 0
rect 510 -13 525 0
<< polycont >>
rect -129 55 -109 75
<< locali >>
rect -100 256 583 260
rect -100 238 -55 256
rect -38 238 0 256
rect 17 238 46 256
rect 63 238 115 256
rect 132 238 170 256
rect 187 238 216 256
rect 233 238 285 256
rect 302 238 340 256
rect 357 238 386 256
rect 403 238 455 256
rect 472 238 510 256
rect 527 238 556 256
rect 573 238 583 256
rect -100 235 583 238
rect -100 234 -40 235
rect 70 234 130 235
rect 240 234 300 235
rect 410 234 470 235
rect -75 218 -40 234
rect 95 218 130 234
rect 265 218 300 234
rect 435 218 470 234
rect -75 210 -5 218
rect -75 207 -30 210
rect -75 189 -69 207
rect -51 189 -30 207
rect -75 188 -30 189
rect -10 188 -5 210
rect -75 168 -5 188
rect -75 165 -30 168
rect -75 147 -69 165
rect -51 147 -30 165
rect -75 146 -30 147
rect -10 146 -5 168
rect -75 126 -5 146
rect -75 123 -30 126
rect -75 105 -69 123
rect -51 105 -30 123
rect -75 104 -30 105
rect -10 104 -5 126
rect -75 96 -5 104
rect 17 210 53 218
rect 17 188 25 210
rect 45 188 53 210
rect 17 168 53 188
rect 17 146 25 168
rect 45 146 53 168
rect 17 126 53 146
rect 17 104 25 126
rect 45 104 53 126
rect 17 96 53 104
rect 95 210 165 218
rect 95 207 140 210
rect 95 189 101 207
rect 119 189 140 207
rect 95 188 140 189
rect 160 188 165 210
rect 95 168 165 188
rect 95 165 140 168
rect 95 147 101 165
rect 119 147 140 165
rect 95 146 140 147
rect 160 146 165 168
rect 95 126 165 146
rect 95 123 140 126
rect 95 105 101 123
rect 119 105 140 123
rect 95 104 140 105
rect 160 104 165 126
rect 95 96 165 104
rect 187 210 223 218
rect 187 188 195 210
rect 215 188 223 210
rect 187 168 223 188
rect 187 146 195 168
rect 215 146 223 168
rect 187 126 223 146
rect 187 104 195 126
rect 215 104 223 126
rect 187 96 223 104
rect 265 210 335 218
rect 265 207 310 210
rect 265 189 271 207
rect 289 189 310 207
rect 265 188 310 189
rect 330 188 335 210
rect 265 168 335 188
rect 265 165 310 168
rect 265 147 271 165
rect 289 147 310 165
rect 265 146 310 147
rect 330 146 335 168
rect 265 126 335 146
rect 265 123 310 126
rect 265 105 271 123
rect 289 105 310 123
rect 265 104 310 105
rect 330 104 335 126
rect 265 96 335 104
rect 357 210 393 218
rect 357 188 365 210
rect 385 188 393 210
rect 357 168 393 188
rect 357 146 365 168
rect 385 146 393 168
rect 357 126 393 146
rect 357 104 365 126
rect 385 104 393 126
rect 357 96 393 104
rect 435 210 505 218
rect 435 207 480 210
rect 435 189 441 207
rect 459 189 480 207
rect 435 188 480 189
rect 500 188 505 210
rect 435 168 505 188
rect 435 165 480 168
rect 435 147 441 165
rect 459 147 480 165
rect 435 146 480 147
rect 500 146 505 168
rect 435 126 505 146
rect 435 123 480 126
rect 435 105 441 123
rect 459 105 480 123
rect 435 104 480 105
rect 500 104 505 126
rect 435 96 505 104
rect 527 210 563 218
rect 527 188 535 210
rect 555 188 563 210
rect 527 168 563 188
rect 527 146 535 168
rect 555 146 563 168
rect 527 126 563 146
rect 527 104 535 126
rect 555 104 563 126
rect 527 96 563 104
rect -137 75 -101 83
rect -137 55 -129 75
rect -109 55 -101 75
rect -137 47 -101 55
rect 24 79 46 96
rect 194 79 216 96
rect 364 79 386 96
rect 534 79 556 96
rect 24 60 556 79
rect 24 40 46 60
rect 194 40 216 60
rect 364 40 386 60
rect 534 40 556 60
rect -75 32 -5 40
rect -75 29 -30 32
rect -75 11 -69 29
rect -51 11 -30 29
rect -75 10 -30 11
rect -10 10 -5 32
rect -75 2 -5 10
rect 17 32 53 40
rect 17 10 25 32
rect 45 10 53 32
rect 17 2 53 10
rect 95 32 165 40
rect 95 29 140 32
rect 95 11 101 29
rect 119 11 140 29
rect 95 10 140 11
rect 160 10 165 32
rect 95 2 165 10
rect 187 32 223 40
rect 187 10 195 32
rect 215 10 223 32
rect 187 2 223 10
rect 265 32 335 40
rect 265 29 310 32
rect 265 11 271 29
rect 289 11 310 29
rect 265 10 310 11
rect 330 10 335 32
rect 265 2 335 10
rect 357 32 393 40
rect 357 10 365 32
rect 385 10 393 32
rect 357 2 393 10
rect 435 32 505 40
rect 435 29 480 32
rect 435 11 441 29
rect 459 11 480 29
rect 435 10 480 11
rect 500 10 505 32
rect 435 2 505 10
rect 527 32 563 40
rect 527 10 535 32
rect 555 10 563 32
rect 527 2 563 10
rect -75 -13 -40 2
rect 95 -13 130 2
rect 265 -13 300 2
rect 435 -13 470 2
rect -100 -15 -40 -13
rect 70 -15 130 -13
rect 240 -15 300 -13
rect 410 -15 470 -13
rect -100 -16 582 -15
rect -100 -34 -55 -16
rect -38 -34 0 -16
rect 17 -34 46 -16
rect 63 -34 115 -16
rect 132 -34 170 -16
rect 187 -34 216 -16
rect 233 -34 285 -16
rect 302 -34 340 -16
rect 357 -34 386 -16
rect 403 -34 455 -16
rect 472 -34 510 -16
rect 527 -34 556 -16
rect 573 -34 582 -16
rect -100 -40 582 -34
<< viali >>
rect -55 238 -38 256
rect 0 238 17 256
rect 46 238 63 256
rect 115 238 132 256
rect 170 238 187 256
rect 216 238 233 256
rect 285 238 302 256
rect 340 238 357 256
rect 386 238 403 256
rect 455 238 472 256
rect 510 238 527 256
rect 556 238 573 256
rect -55 -34 -38 -16
rect 0 -34 17 -16
rect 46 -34 63 -16
rect 115 -34 132 -16
rect 170 -34 187 -16
rect 216 -34 233 -16
rect 285 -34 302 -16
rect 340 -34 357 -16
rect 386 -34 403 -16
rect 455 -34 472 -16
rect 510 -34 527 -16
rect 556 -34 573 -16
<< metal1 >>
rect -100 256 583 260
rect -100 238 -55 256
rect -38 238 0 256
rect 17 238 46 256
rect 63 238 115 256
rect 132 238 170 256
rect 187 238 216 256
rect 233 238 285 256
rect 302 238 340 256
rect 357 238 386 256
rect 403 238 455 256
rect 472 238 510 256
rect 527 238 556 256
rect 573 238 583 256
rect -100 234 583 238
rect -100 -16 583 -13
rect -100 -34 -55 -16
rect -38 -34 0 -16
rect 17 -34 46 -16
rect 63 -34 115 -16
rect 132 -34 170 -16
rect 187 -34 216 -16
rect 233 -34 285 -16
rect 302 -34 340 -16
rect 357 -34 386 -16
rect 403 -34 455 -16
rect 472 -34 510 -16
rect 527 -34 556 -16
rect 573 -34 583 -16
rect -100 -40 583 -34
<< labels >>
rlabel metal1 -99 247 -99 247 1 vdd
port 1 n
rlabel metal1 -99 -27 -99 -27 1 vss
port 2 n
rlabel locali -136 65 -136 65 3 in
port 3 e
rlabel locali 555 69 555 69 1 out
port 4 n
<< end >>
